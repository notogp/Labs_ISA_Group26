library verilog;
use verilog.vl_types.all;
entity tb_fir_unfolded is
end tb_fir_unfolded;
